module upsample_test;
  integer  satId,i;
  real sample_count;
  real sampling_freq = 18548387;
  real code_length = 10230;
  real code_freq_basis = 1023000;
  real ind_array[];
  initial begin
    sample_count = sampling_freq/(code_freq_basis/code_length);
    ind_array = new[sample_count];
    for (i=0; i<sample_count; i=i+1) begin
      //ind_array[i] = int'((i*code_freq_basis)/sampling_freq);
      ind_array[i] = $rtoi((i*code_freq_basis)/sampling_freq);
    end
    //$display("index_val = %g",ind_array[91]);
    for(int i=0; i< 100;i=i+1) begin
      $write("%g,",ind_array[i]); 
      //$write("\n"); 
    end
    $display("sample_count = %g",sample_count);
  end
endmodule
