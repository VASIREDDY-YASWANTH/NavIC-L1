
`define pi 16'b011_0010010000111
module Cosin
  #(parameter DEPTH=256,parameter WIDTH = 16);

//bit signed [WIDTH-1:0] array[DEPTH] = '{16'b0_000000000000000, 16'b0_000110010001011, 16'b0_001100011111001, 16'b0_010010100101000, 16'b0_011000011111100, 16'b0_011110001010110, 16'b0_100011100011101, 16'b0_101000100110100, 16'b0_101101010000010, 16'b0_110001011110001, 16'b0_110101001101110, 16'b0_111000011100010, 16'b0_111011001000010, 16'b0_111101001111011, 16'b0_111110110001010, 16'b0_111111101100010};
bit signed [WIDTH-1:0] array[DEPTH] = '{16'b0_000000000000000,                               
16'b0_000000011001001,                              
16'b0_000000110010010,                               
16'b0_000001001011011,                               
16'b0_000001100100100,                               
16'b0_000001111101101,                               
16'b0_000010010110110,                               
16'b0_000010101111111,                               
16'b0_000011001000111,                               
16'b0_000011100010000,                               
16'b0_000011111011001,                               
16'b0_000100010100010,                               
16'b0_000100101101010,                               
16'b0_000101000110011,                               
16'b0_000101011111011,                               
16'b0_000101111000011,                               
16'b0_000110010001011,                               
16'b0_000110101010011,                               
16'b0_000111000011011,                               
16'b0_000111011100011,                               
16'b0_000111110101011,                               
16'b0_001000001110010,                               
16'b0_001000100111001,                               
16'b0_001001000000001,                               
16'b0_001001011001000,                               
16'b0_001001110001110,                               
16'b0_001010001010101,                               
16'b0_001010100011011,                               
16'b0_001010111100010,                               
16'b0_001011010101000,                               
16'b0_001011101101101,                               
16'b0_001100000110011,                               
16'b0_001100011111000,                               
16'b0_001100110111101,                               
16'b0_001101010000010,                               
16'b0_001101101000111,                               
16'b0_001110000001011,                               
16'b0_001110011001111,                               
16'b0_001110110010011,                               
16'b0_001111001010110,                               
16'b0_001111100011001,                               
16'b0_001111111011100,                               
16'b0_010000010011111,                               
16'b0_010000101100001,                               
16'b0_010001000100011,                               
16'b0_010001011100101,                               
16'b0_010001110100110,                               
16'b0_010010001100111,                               
16'b0_010010100101000,                               
16'b0_010010111101000,                               
16'b0_010011010101000,                               
16'b0_010011101100111,                               
16'b0_010100000100110,                               
16'b0_010100011100101,                               
16'b0_010100110100011,                               
16'b0_010101001100001,                               
16'b0_010101100011111,                               
16'b0_010101111011100,                               
16'b0_010110010011000,                               
16'b0_010110101010101,                               
16'b0_010111000010001,                               
16'b0_010111011001100,                               
16'b0_010111110000111,                               
16'b0_011000001000001,                               
16'b0_011000011111011,                               
16'b0_011000110110101,                               
16'b0_011001001101110,                               
16'b0_011001100100110,                               
16'b0_011001111011110,                               
16'b0_011010010010110,                               
16'b0_011010101001101,                               
16'b0_011011000000100,                               
16'b0_011011010111010,                               
16'b0_011011101101111,                               
16'b0_011100000100100,                               
16'b0_011100011011000,                               
16'b0_011100110001100,                               
16'b0_011101001000000,                               
16'b0_011101011110010,                               
16'b0_011101110100101,                               
16'b0_011110001010110,                               
16'b0_011110100000111,                               
16'b0_011110110111000,                               
16'b0_011111001101000,                               
16'b0_011111100010111,                               
16'b0_011111111000101,                               
16'b0_100000001110011,                               
16'b0_100000100100001,                               
16'b0_100000111001110,                               
16'b0_100001001111010,                               
16'b0_100001100100101,                               
16'b0_100001111010000,                               
16'b0_100010001111010,                               
16'b0_100010100100100,                               
16'b0_100010111001101,                               
16'b0_100011001110101,                               
16'b0_100011100011100,                               
16'b0_100011111000011,                               
16'b0_100100001101001,                               
16'b0_100100100001111,                               
16'b0_100100110110100,                               
16'b0_100101001011000,                               
16'b0_100101011111011,                               
16'b0_100101110011110,                               
16'b0_100110000111111,                               
16'b0_100110011100001,                               
16'b0_100110110000001,                               
16'b0_100111000100001,                               
16'b0_100111010111111,                               
16'b0_100111101011110,                               
16'b0_100111111111011,                               
16'b0_101000010010111,                               
16'b0_101000100110011,                               
16'b0_101000111001110,                               
16'b0_101001001101001,                               
16'b0_101001100000010,                               
16'b0_101001110011011,                               
16'b0_101010000110011,                               
16'b0_101010011001010,                               
16'b0_101010101100000,                               
16'b0_101010111110101,                               
16'b0_101011010001010,                               
16'b0_101011100011101,                               
16'b0_101011110110000,                               
16'b0_101100001000010,                               
16'b0_101100011010100,                               
16'b0_101100101100100,                               
16'b0_101100111110011,                               
16'b0_101101010000010,                               
16'b0_101101100010000,                               
16'b0_101101110011101,                               
16'b0_101110000101001,                               
16'b0_101110010110100,                               
16'b0_101110100111110,                               
16'b0_101110111000111,                               
16'b0_101111001010000,                               
16'b0_101111011010111,                               
16'b0_101111101011110,                               
16'b0_101111111100011,                               
16'b0_110000001101000,                               
16'b0_110000011101100,                               
16'b0_110000101101111,                               
16'b0_110000111110001,                               
16'b0_110001001110001,                               
16'b0_110001011110010,                               
16'b0_110001101110001,                               
16'b0_110001111101111,                               
16'b0_110010001101100,                               
16'b0_110010011101000,                               
16'b0_110010101100011,                               
16'b0_110010111011101,                               
16'b0_110011001010111,                               
16'b0_110011011001111,                               
16'b0_110011101000110,                               
16'b0_110011110111101,                               
16'b0_110100000110010,                               
16'b0_110100010100110,                               
16'b0_110100100011001,                               
16'b0_110100110001100,                               
16'b0_110100111111101,                               
16'b0_110101001101101,                               
16'b0_110101011011100,                               
16'b0_110101101001010,                               
16'b0_110101110111000,                               
16'b0_110110000100100,                               
16'b0_110110010001111,                               
16'b0_110110011111001,                               
16'b0_110110101100010,                               
16'b0_110110111001010,                               
16'b0_110111000110000,                               
16'b0_110111010010110,                               
16'b0_110111011111011,                               
16'b0_110111101011111,                               
16'b0_110111111000001,                               
16'b0_111000000100011,                               
16'b0_111000010000011,                               
16'b0_111000011100010,                               
16'b0_111000101000001,                               
16'b0_111000110011110,                               
16'b0_111000111111010,                               
16'b0_111001001010101,                               
16'b0_111001010101111,                               
16'b0_111001100000111,                               
16'b0_111001101011111,                               
16'b0_111001110110101,                               
16'b0_111010000001011,                               
16'b0_111010001011111,                               
16'b0_111010010110010,                               
16'b0_111010100000100,                               
16'b0_111010101010101,                               
16'b0_111010110100101,                               
16'b0_111010111110100,                               
16'b0_111011001000001,                               
16'b0_111011010001110,                               
16'b0_111011011011001,                               
16'b0_111011100100011,                               
16'b0_111011101101100,                               
16'b0_111011110110100,                               
16'b0_111011111111010,                               
16'b0_111100001000000,                               
16'b0_111100010000100,                               
16'b0_111100011000111,                               
16'b0_111100100001001,                               
16'b0_111100101001010,                               
16'b0_111100110001010,                               
16'b0_111100111001000,                               
16'b0_111101000000101,                               
16'b0_111101001000010,                               
16'b0_111101001111101,                               
16'b0_111101010110110,                               
16'b0_111101011101111,                               
16'b0_111101100100110,                               
16'b0_111101101011101,                               
16'b0_111101110010010,                               
16'b0_111101111000101,                               
16'b0_111101111111000,                               
16'b0_111110000101001,                               
16'b0_111110001011010,                               
16'b0_111110010001001,                               
16'b0_111110010110111,                               
16'b0_111110011100011,                               
16'b0_111110100001111,                               
16'b0_111110100111001,                               
16'b0_111110101100010,                               
16'b0_111110110001010,                               
16'b0_111110110110000,                               
16'b0_111110111010110,                               
16'b0_111110111111010,                               
16'b0_111111000011101,                               
16'b0_111111000111111,                               
16'b0_111111001011111,                               
16'b0_111111001111111,                               
16'b0_111111010011101,                               
16'b0_111111010111010,                               
16'b0_111111011010101,                               
16'b0_111111011110000,                               
16'b0_111111100001001,                               
16'b0_111111100100001,                               
16'b0_111111100111000,                               
16'b0_111111101001101,                               
16'b0_111111101100010,                               
16'b0_111111101110101,                               
16'b0_111111110000111,                               
16'b0_111111110010111,                               
16'b0_111111110100111,                               
16'b0_111111110110101,                               
16'b0_111111111000010,                               
16'b0_111111111001110,                               
16'b0_111111111011000,                               
16'b0_111111111100001,                               
16'b0_111111111101001,                               
16'b0_111111111110000,                               
16'b0_111111111110110,                               
16'b0_111111111111010,                               
16'b0_111111111111101,                               
16'b1_000000000000000                               
};
   
localparam SF = 2.0**-15.0;
localparam SF1 = 2.0**-13.0;
int n = 1;
// function for Sine Computation
  function bit signed [WIDTH-1:0] sin_tab;
	input bit [31:0] angle; 
	int index,x1,x2;
	real indexr,x;
	bit signed [WIDTH-1:0] y1,y2,y;
    
    begin
      // changing angle value in the range of {0 to pi/2}
      while (angle>(2*`pi))begin
        angle = angle-(2*`pi);
      end
      $display("angle=%g",angle*SF1);
      //finding corresponding index for given angle 
      index = int'(angle/(`pi/(2*DEPTH)));
      indexr = $itor(angle*SF1)/($itor(`pi*SF1)/(2*DEPTH)) ;
      index= $floor(indexr);
      x=indexr-index;
      $display("Index = %0d",index);
      //finding index lies in which Quadrant
      if (index<DEPTH)begin             //1st Quadrant
        $display("Index = %0d",index);
        sin_tab = array[index];
      end
      else if ((2*DEPTH)>index)begin    //2nd Quadrant
        index = ((2*DEPTH)-1)-index;
	x=1-x;
        $display("Index = %0d",index);
        sin_tab = array[index];
      end
      else if ((3*DEPTH)>index)begin    //3rd Quadrant
        index = index-(2*DEPTH);
        $display("Index = %0d",index);
        sin_tab = -array[index];
      end
      else if ((4*DEPTH)>index)begin     //4th Quadrant
        index = ((4*DEPTH)-1)-index;
	x=1-x;
        $display("Index = %0d",index);
        sin_tab = -array[index];
      end

$display("Indexr = %0f",indexr);
$display("x = %0f", x );
x1=index;
x2=index+1;

if (x1<DEPTH)begin
        y1 = array[x1];
      end
      else if ((2*DEPTH)>x1)begin
        x1 = ((2*DEPTH)-1)-x1;
        y1 = array[x1];
      end
      else if ((3*DEPTH)>x1)begin
        x1 = x1-(2*DEPTH);
        y1 = -array[x1];
      end
      else if ((4*DEPTH)>x1)begin
        x1 = ((4*DEPTH)-1)-x1;
        y1 = -array[x1];
      end

if (x2<DEPTH)begin
        y2 = array[x2];
      end
      else if ((2*DEPTH)>x2)begin
        x2 = ((2*DEPTH)-1)-x2;
        y2 = array[x2];
      end
      else if ((3*DEPTH)>x2)begin
        x2 = x2-(2*DEPTH);
        y2 = -array[x2];
      end
      else if ((4*DEPTH)>x2)begin
        x2 = ((4*DEPTH)-1)-x2;
        y2 = -array[x2];
      end

//Interpolation
$display("x2,y2 = %0d, %0f ",x2,y2*SF);
$display("x1,y1 = %0d, %0f ",x1,y1*SF);
y=y1+(y2-y1)*x;
$display("y = %0f",y*SF);

    end
  endfunction

//function for Cosine Computation
  function bit signed [WIDTH-1:0] cos_tab;
    input bit [15:0] angle_1;
    begin
      cos_tab = sin_tab(angle_1+(`pi/2));
    end
  endfunction

// Main Function
  initial begin
    bit [31:0] val;
    bit signed [15:0] result1,result2;
	//for(int i=2;i<16;i++)begin
     val = ((`pi)/13);
    //$display("val=%g",val*SF1);
	
    result1 = sin_tab(val);
   // $display("sin(%0f) = %0b", val*SF1, result1);
    $display("sin(%0f) = %0g\n  %f", val*SF1, result1*SF,$itor(result1*SF) - $sin(val));
   // result2 = cos_tab(val);
    //$display("cos(%0f) = %0b", val*SF1, result2);
   // $display("cos(%0f) = %0g", val*SF1, result2*SF);
  
  end
endmodule